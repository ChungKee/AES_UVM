interface AES_interface;
    logic clk;
    logic rst;
    logic [127:0]P;
    logic [127:0]K;
    logic [127:0]C;
    logic valid;
endinterface
